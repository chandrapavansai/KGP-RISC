`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:17:17 10/08/2021 
// Design Name: 
// Module Name:    mux_2_1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
//
// Assignment 6
// Semester no 5
// Group No 51
// Question no 1
// KPSM Surya
// Pavan Sai Chandra
//
//////////////////////////////////////////////////////////////////////////////////
module mux_2_1(
    input sel,
    input A,
    input B,
    output o
    );
	 assign o = (sel)? A: B;

endmodule
